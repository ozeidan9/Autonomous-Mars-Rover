// Qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module Qsys (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //      alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                                 .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                                 .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                                 .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                                 .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                                 .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                                 .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                                 .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                                 .vid_v
		input  wire        altpll_0_areset_conduit_export,            //          altpll_0_areset_conduit.export
		output wire        altpll_0_locked_conduit_export,            //          altpll_0_locked_conduit.export
		input  wire        clk_clk,                                   //                              clk.clk
		output wire        clk_sdram_clk,                             //                        clk_sdram.clk
		output wire        clk_vga_clk,                               //                          clk_vga.clk
		output wire        d8m_xclkin_clk,                            //                       d8m_xclkin.clk
		output wire [15:0] eee_imgproc_0_avalon_slave_0_readdata,     //     eee_imgproc_0_avalon_slave_0.readdata
		input  wire        eee_imgproc_0_conduit_mode_new_signal,     //       eee_imgproc_0_conduit_mode.new_signal
		input  wire [15:0] eee_imgproc_0_conduit_mode_new_signal_1,   //                                 .new_signal_1
		inout  wire        i2c_opencores_camera_export_scl_pad_io,    //      i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,    //                                 .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,      //        i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,      //                                 .sda_pad_io
		input  wire [1:0]  key_external_connection_export,            //          key_external_connection.export
		output wire [9:0]  led_external_connection_export,            //          led_external_connection.export
		output wire        mipi_pwdn_n_external_connection_export,    //  mipi_pwdn_n_external_connection.export
		output wire        mipi_reset_n_external_connection_export,   // mipi_reset_n_external_connection.export
		input  wire        reset_reset_n,                             //                            reset.reset_n
		output wire [12:0] sdram_wire_addr,                           //                       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                                 .ba
		output wire        sdram_wire_cas_n,                          //                                 .cas_n
		output wire        sdram_wire_cke,                            //                                 .cke
		output wire        sdram_wire_cs_n,                           //                                 .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                                 .dq
		output wire [1:0]  sdram_wire_dqm,                            //                                 .dqm
		output wire        sdram_wire_ras_n,                          //                                 .ras_n
		output wire        sdram_wire_we_n,                           //                                 .we_n
		input  wire [9:0]  sw_external_connection_export,             //           sw_external_connection.export
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_sda,  //     terasic_auto_focus_0_conduit.vcm_i2c_sda
		input  wire        terasic_auto_focus_0_conduit_clk50,        //                                 .clk50
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_scl,  //                                 .vcm_i2c_scl
		input  wire [11:0] terasic_camera_0_conduit_end_D,            //     terasic_camera_0_conduit_end.D
		input  wire        terasic_camera_0_conduit_end_FVAL,         //                                 .FVAL
		input  wire        terasic_camera_0_conduit_end_LVAL,         //                                 .LVAL
		input  wire        terasic_camera_0_conduit_end_PIXCLK,       //                                 .PIXCLK
		input  wire        uart_0_rx_tx_rxd,                          //                     uart_0_rx_tx.rxd
		output wire        uart_0_rx_tx_txd                           //                                 .txd
	);

	wire         terasic_camera_0_avalon_streaming_source_valid;                    // TERASIC_CAMERA_0:st_valid -> alt_vip_vfb_0:din_valid
	wire  [23:0] terasic_camera_0_avalon_streaming_source_data;                     // TERASIC_CAMERA_0:st_data -> alt_vip_vfb_0:din_data
	wire         terasic_camera_0_avalon_streaming_source_ready;                    // alt_vip_vfb_0:din_ready -> TERASIC_CAMERA_0:st_ready
	wire         terasic_camera_0_avalon_streaming_source_startofpacket;            // TERASIC_CAMERA_0:st_sop -> alt_vip_vfb_0:din_startofpacket
	wire         terasic_camera_0_avalon_streaming_source_endofpacket;              // TERASIC_CAMERA_0:st_eop -> alt_vip_vfb_0:din_endofpacket
	wire         eee_imgproc_0_avalon_streaming_source_valid;                       // EEE_IMGPROC_0:source_valid -> alt_vip_itc_0:is_valid
	wire  [23:0] eee_imgproc_0_avalon_streaming_source_data;                        // EEE_IMGPROC_0:source_data -> alt_vip_itc_0:is_data
	wire         eee_imgproc_0_avalon_streaming_source_ready;                       // alt_vip_itc_0:is_ready -> EEE_IMGPROC_0:source_ready
	wire         eee_imgproc_0_avalon_streaming_source_startofpacket;               // EEE_IMGPROC_0:source_sop -> alt_vip_itc_0:is_sop
	wire         eee_imgproc_0_avalon_streaming_source_endofpacket;                 // EEE_IMGPROC_0:source_eop -> alt_vip_itc_0:is_eop
	wire         terasic_auto_focus_0_dout_valid;                                   // TERASIC_AUTO_FOCUS_0:source_valid -> EEE_IMGPROC_0:sink_valid
	wire  [23:0] terasic_auto_focus_0_dout_data;                                    // TERASIC_AUTO_FOCUS_0:source_data -> EEE_IMGPROC_0:sink_data
	wire         terasic_auto_focus_0_dout_ready;                                   // EEE_IMGPROC_0:sink_ready -> TERASIC_AUTO_FOCUS_0:source_ready
	wire         terasic_auto_focus_0_dout_startofpacket;                           // TERASIC_AUTO_FOCUS_0:source_sop -> EEE_IMGPROC_0:sink_sop
	wire         terasic_auto_focus_0_dout_endofpacket;                             // TERASIC_AUTO_FOCUS_0:source_eop -> EEE_IMGPROC_0:sink_eop
	wire         alt_vip_vfb_0_dout_valid;                                          // alt_vip_vfb_0:dout_valid -> TERASIC_AUTO_FOCUS_0:sink_valid
	wire  [23:0] alt_vip_vfb_0_dout_data;                                           // alt_vip_vfb_0:dout_data -> TERASIC_AUTO_FOCUS_0:sink_data
	wire         alt_vip_vfb_0_dout_ready;                                          // TERASIC_AUTO_FOCUS_0:sink_ready -> alt_vip_vfb_0:dout_ready
	wire         alt_vip_vfb_0_dout_startofpacket;                                  // alt_vip_vfb_0:dout_startofpacket -> TERASIC_AUTO_FOCUS_0:sink_sop
	wire         alt_vip_vfb_0_dout_endofpacket;                                    // alt_vip_vfb_0:dout_endofpacket -> TERASIC_AUTO_FOCUS_0:sink_eop
	wire         altpll_0_c2_clk;                                                   // altpll_0:c2 -> [EEE_IMGPROC_0:clk, TERASIC_AUTO_FOCUS_0:clk, TERASIC_CAMERA_0:clk, alt_vip_itc_0:is_clk, alt_vip_vfb_0:clock, mm_interconnect_0:altpll_0_c2_clk, mm_interconnect_1:altpll_0_c2_clk, rst_controller:clk, sdram:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                                   // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                                // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                                // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [18:0] nios2_gen2_data_master_address;                                    // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                 // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                       // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                              // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                      // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                  // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                            // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [18:0] nios2_gen2_instruction_master_address;                             // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                                // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect;    // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata;      // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest;   // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address;       // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write;         // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata;     // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect;  // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata;    // i2c_opencores_camera:wb_dat_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest; // i2c_opencores_camera:wb_ack_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address;     // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write;       // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata;   // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;               // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;             // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;          // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;              // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                 // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;            // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect;         // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect -> TERASIC_AUTO_FOCUS_0:s_chipselect
	wire  [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata;           // TERASIC_AUTO_FOCUS_0:s_readdata -> mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata
	wire   [2:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address;            // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_address -> TERASIC_AUTO_FOCUS_0:s_address
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read;               // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_read -> TERASIC_AUTO_FOCUS_0:s_read
	wire         mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write;              // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_write -> TERASIC_AUTO_FOCUS_0:s_write
	wire  [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata;          // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata -> TERASIC_AUTO_FOCUS_0:s_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                     // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                      // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                         // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                        // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                    // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                             // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                               // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                  // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                              // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                               // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                 // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                  // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                    // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                  // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                   // mm_interconnect_0:sw_s1_address -> sw:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                 // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                  // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_mipi_reset_n_s1_chipselect;                      // mm_interconnect_0:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_readdata;                        // mipi_reset_n:readdata -> mm_interconnect_0:mipi_reset_n_s1_readdata
	wire   [1:0] mm_interconnect_0_mipi_reset_n_s1_address;                         // mm_interconnect_0:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire         mm_interconnect_0_mipi_reset_n_s1_write;                           // mm_interconnect_0:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire  [31:0] mm_interconnect_0_mipi_reset_n_s1_writedata;                       // mm_interconnect_0:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire         mm_interconnect_0_mipi_pwdn_n_s1_chipselect;                       // mm_interconnect_0:mipi_pwdn_n_s1_chipselect -> mipi_pwdn_n:chipselect
	wire  [31:0] mm_interconnect_0_mipi_pwdn_n_s1_readdata;                         // mipi_pwdn_n:readdata -> mm_interconnect_0:mipi_pwdn_n_s1_readdata
	wire   [1:0] mm_interconnect_0_mipi_pwdn_n_s1_address;                          // mm_interconnect_0:mipi_pwdn_n_s1_address -> mipi_pwdn_n:address
	wire         mm_interconnect_0_mipi_pwdn_n_s1_write;                            // mm_interconnect_0:mipi_pwdn_n_s1_write -> mipi_pwdn_n:write_n
	wire  [31:0] mm_interconnect_0_mipi_pwdn_n_s1_writedata;                        // mm_interconnect_0:mipi_pwdn_n_s1_writedata -> mipi_pwdn_n:writedata
	wire         mm_interconnect_0_eee_imgproc_0_s1_chipselect;                     // mm_interconnect_0:EEE_IMGPROC_0_s1_chipselect -> EEE_IMGPROC_0:s_chipselect
	wire  [31:0] mm_interconnect_0_eee_imgproc_0_s1_readdata;                       // EEE_IMGPROC_0:s_readdata -> mm_interconnect_0:EEE_IMGPROC_0_s1_readdata
	wire   [2:0] mm_interconnect_0_eee_imgproc_0_s1_address;                        // mm_interconnect_0:EEE_IMGPROC_0_s1_address -> EEE_IMGPROC_0:s_address
	wire         mm_interconnect_0_eee_imgproc_0_s1_read;                           // mm_interconnect_0:EEE_IMGPROC_0_s1_read -> EEE_IMGPROC_0:s_read
	wire         mm_interconnect_0_eee_imgproc_0_s1_write;                          // mm_interconnect_0:EEE_IMGPROC_0_s1_write -> EEE_IMGPROC_0:s_write
	wire  [31:0] mm_interconnect_0_eee_imgproc_0_s1_writedata;                      // mm_interconnect_0:EEE_IMGPROC_0_s1_writedata -> EEE_IMGPROC_0:s_writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                            // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                              // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                               // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                  // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                         // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                 // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                             // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         alt_vip_vfb_0_read_master_waitrequest;                             // mm_interconnect_1:alt_vip_vfb_0_read_master_waitrequest -> alt_vip_vfb_0:read_master_av_waitrequest
	wire  [31:0] alt_vip_vfb_0_read_master_readdata;                                // mm_interconnect_1:alt_vip_vfb_0_read_master_readdata -> alt_vip_vfb_0:read_master_av_readdata
	wire  [31:0] alt_vip_vfb_0_read_master_address;                                 // alt_vip_vfb_0:read_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_read_master_address
	wire         alt_vip_vfb_0_read_master_read;                                    // alt_vip_vfb_0:read_master_av_read -> mm_interconnect_1:alt_vip_vfb_0_read_master_read
	wire         alt_vip_vfb_0_read_master_readdatavalid;                           // mm_interconnect_1:alt_vip_vfb_0_read_master_readdatavalid -> alt_vip_vfb_0:read_master_av_readdatavalid
	wire   [2:0] alt_vip_vfb_0_read_master_burstcount;                              // alt_vip_vfb_0:read_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_read_master_burstcount
	wire         alt_vip_vfb_0_write_master_waitrequest;                            // mm_interconnect_1:alt_vip_vfb_0_write_master_waitrequest -> alt_vip_vfb_0:write_master_av_waitrequest
	wire  [31:0] alt_vip_vfb_0_write_master_address;                                // alt_vip_vfb_0:write_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_write_master_address
	wire         alt_vip_vfb_0_write_master_write;                                  // alt_vip_vfb_0:write_master_av_write -> mm_interconnect_1:alt_vip_vfb_0_write_master_write
	wire  [31:0] alt_vip_vfb_0_write_master_writedata;                              // alt_vip_vfb_0:write_master_av_writedata -> mm_interconnect_1:alt_vip_vfb_0_write_master_writedata
	wire   [2:0] alt_vip_vfb_0_write_master_burstcount;                             // alt_vip_vfb_0:write_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_write_master_burstcount
	wire         mm_interconnect_1_sdram_s1_chipselect;                             // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_1_sdram_s1_readdata;                               // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire         mm_interconnect_1_sdram_s1_waitrequest;                            // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_1_sdram_s1_address;                                // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_1_sdram_s1_read;                                   // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_1_sdram_s1_byteenable;                             // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                          // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire         mm_interconnect_1_sdram_s1_write;                                  // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_1_sdram_s1_writedata;                              // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire         irq_mapper_receiver0_irq;                                          // i2c_opencores_mipi:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // i2c_opencores_camera:wb_inta_o -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                          // timer:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                          // uart_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_irq_irq;                                                // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [EEE_IMGPROC_0:reset_n, TERASIC_AUTO_FOCUS_0:reset_n, TERASIC_CAMERA_0:reset_n, alt_vip_itc_0:rst, alt_vip_vfb_0:reset, mm_interconnect_0:TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_vfb_0_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         nios2_gen2_debug_reset_request_reset;                              // nios2_gen2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [i2c_opencores_camera:wb_rst_i, i2c_opencores_mipi:wb_rst_i, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, led:reset_n, mipi_pwdn_n:reset_n, mipi_reset_n:reset_n, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sw:reset_n, sysid_qsys:reset_n, timer:reset_n, uart_0:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                            // rst_controller_002:reset_req -> [nios2_gen2:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	EEE_IMGPROC #(
		.IMAGE_W         (13'b0001010000000),
		.IMAGE_H         (13'b0000111100000),
		.MESSAGE_BUF_MAX (256),
		.MSG_INTERVAL    (6),
		.BB_COL_DEFAULT  (26'b00000000001111111100000000)
	) eee_imgproc_0 (
		.clk                (altpll_0_c2_clk),                                     //                   clock.clk
		.reset_n            (~rst_controller_reset_out_reset),                     //                   reset.reset_n
		.sink_data          (terasic_auto_focus_0_dout_data),                      //   avalon_streaming_sink.data
		.sink_valid         (terasic_auto_focus_0_dout_valid),                     //                        .valid
		.sink_ready         (terasic_auto_focus_0_dout_ready),                     //                        .ready
		.sink_sop           (terasic_auto_focus_0_dout_startofpacket),             //                        .startofpacket
		.sink_eop           (terasic_auto_focus_0_dout_endofpacket),               //                        .endofpacket
		.source_data        (eee_imgproc_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.source_eop         (eee_imgproc_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.source_ready       (eee_imgproc_0_avalon_streaming_source_ready),         //                        .ready
		.source_sop         (eee_imgproc_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.source_valid       (eee_imgproc_0_avalon_streaming_source_valid),         //                        .valid
		.s_chipselect       (mm_interconnect_0_eee_imgproc_0_s1_chipselect),       //                      s1.chipselect
		.s_read             (mm_interconnect_0_eee_imgproc_0_s1_read),             //                        .read
		.s_write            (mm_interconnect_0_eee_imgproc_0_s1_write),            //                        .write
		.s_readdata         (mm_interconnect_0_eee_imgproc_0_s1_readdata),         //                        .readdata
		.s_writedata        (mm_interconnect_0_eee_imgproc_0_s1_writedata),        //                        .writedata
		.s_address          (mm_interconnect_0_eee_imgproc_0_s1_address),          //                        .address
		.mode               (eee_imgproc_0_conduit_mode_new_signal),               //            conduit_mode.new_signal
		.byte_data_received (eee_imgproc_0_conduit_mode_new_signal_1),             //                        .new_signal_1
		.outbuffer          (eee_imgproc_0_avalon_slave_0_readdata)                //          avalon_slave_0.readdata
	);

	TERASIC_AUTO_FOCUS #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_auto_focus_0 (
		.clk          (altpll_0_c2_clk),                                           //   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                           //   reset.reset_n
		.s_chipselect (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect), // mm_ctrl.chipselect
		.s_read       (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),       //        .read
		.s_write      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),      //        .write
		.s_readdata   (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),   //        .readdata
		.s_writedata  (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),  //        .writedata
		.s_address    (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),    //        .address
		.sink_data    (alt_vip_vfb_0_dout_data),                                   //     din.data
		.sink_valid   (alt_vip_vfb_0_dout_valid),                                  //        .valid
		.sink_ready   (alt_vip_vfb_0_dout_ready),                                  //        .ready
		.sink_sop     (alt_vip_vfb_0_dout_startofpacket),                          //        .startofpacket
		.sink_eop     (alt_vip_vfb_0_dout_endofpacket),                            //        .endofpacket
		.source_data  (terasic_auto_focus_0_dout_data),                            //    dout.data
		.source_valid (terasic_auto_focus_0_dout_valid),                           //        .valid
		.source_ready (terasic_auto_focus_0_dout_ready),                           //        .ready
		.source_sop   (terasic_auto_focus_0_dout_startofpacket),                   //        .startofpacket
		.source_eop   (terasic_auto_focus_0_dout_endofpacket),                     //        .endofpacket
		.vcm_i2c_sda  (terasic_auto_focus_0_conduit_vcm_i2c_sda),                  // Conduit.vcm_i2c_sda
		.clk50        (terasic_auto_focus_0_conduit_clk50),                        //        .clk50
		.vcm_i2c_scl  (terasic_auto_focus_0_conduit_vcm_i2c_scl)                   //        .vcm_i2c_scl
	);

	TERASIC_CAMERA #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_camera_0 (
		.clk           (altpll_0_c2_clk),                                        //             clock_reset.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //       clock_reset_reset.reset_n
		.CAMERA_D      (terasic_camera_0_conduit_end_D),                         //             conduit_end.export
		.CAMERA_FVAL   (terasic_camera_0_conduit_end_FVAL),                      //                        .export
		.CAMERA_LVAL   (terasic_camera_0_conduit_end_LVAL),                      //                        .export
		.CAMERA_PIXCLK (terasic_camera_0_conduit_end_PIXCLK),                    //                        .export
		.st_data       (terasic_camera_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.st_sop        (terasic_camera_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.st_eop        (terasic_camera_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.st_ready      (terasic_camera_0_avalon_streaming_source_ready),         //                        .ready
		.st_valid      (terasic_camera_0_avalon_streaming_source_valid)          //                        .valid
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (640),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (639),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (10),
		.V_BACK_PORCH                  (33),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (altpll_0_c2_clk),                                     //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),                      // is_clk_rst_reset.reset
		.is_data       (eee_imgproc_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (eee_imgproc_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (eee_imgproc_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (eee_imgproc_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (eee_imgproc_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                 //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),               //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),           //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),              //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),              //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                   //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                   //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                    //                 .export
	);

	Qsys_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (altpll_0_c2_clk),                                        //        clock.clk
		.reset                        (rst_controller_reset_out_reset),                         //        reset.reset
		.din_ready                    (terasic_camera_0_avalon_streaming_source_ready),         //          din.ready
		.din_valid                    (terasic_camera_0_avalon_streaming_source_valid),         //             .valid
		.din_data                     (terasic_camera_0_avalon_streaming_source_data),          //             .data
		.din_startofpacket            (terasic_camera_0_avalon_streaming_source_startofpacket), //             .startofpacket
		.din_endofpacket              (terasic_camera_0_avalon_streaming_source_endofpacket),   //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),                               //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),                               //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),                                //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),                       //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),                         //             .endofpacket
		.read_master_av_address       (alt_vip_vfb_0_read_master_address),                      //  read_master.address
		.read_master_av_read          (alt_vip_vfb_0_read_master_read),                         //             .read
		.read_master_av_waitrequest   (alt_vip_vfb_0_read_master_waitrequest),                  //             .waitrequest
		.read_master_av_readdatavalid (alt_vip_vfb_0_read_master_readdatavalid),                //             .readdatavalid
		.read_master_av_readdata      (alt_vip_vfb_0_read_master_readdata),                     //             .readdata
		.read_master_av_burstcount    (alt_vip_vfb_0_read_master_burstcount),                   //             .burstcount
		.write_master_av_address      (alt_vip_vfb_0_write_master_address),                     // write_master.address
		.write_master_av_write        (alt_vip_vfb_0_write_master_write),                       //             .write
		.write_master_av_writedata    (alt_vip_vfb_0_write_master_writedata),                   //             .writedata
		.write_master_av_waitrequest  (alt_vip_vfb_0_write_master_waitrequest),                 //             .waitrequest
		.write_master_av_burstcount   (alt_vip_vfb_0_write_master_burstcount)                   //             .burstcount
	);

	Qsys_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (),                                               //                    c0.clk
		.c1                 (clk_sdram_clk),                                  //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.c3                 (clk_vga_clk),                                    //                    c3.clk
		.c4                 (d8m_xclkin_clk),                                 //                    c4.clk
		.areset             (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_0_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (clk_clk),                                                           //            clock.clk
		.wb_rst_i   (rst_controller_002_reset_out_reset),                                //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver1_irq)                                           // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (clk_clk),                                                         //            clock.clk
		.wb_rst_i   (rst_controller_002_reset_out_reset),                              //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                         // interrupt_sender.irq
	);

	Qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	Qsys_key key (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	Qsys_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	Qsys_mipi_pwdn_n mipi_pwdn_n (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mipi_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_pwdn_n_external_connection_export)       // external_connection.export
	);

	Qsys_mipi_pwdn_n mipi_reset_n (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	Qsys_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	Qsys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	Qsys_sdram sdram (
		.clk            (altpll_0_c2_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Qsys_sw sw (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_external_connection_export)        // external_connection.export
	);

	Qsys_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	Qsys_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	Qsys_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_rx_tx_rxd),                          // external_connection.export
		.txd           (uart_0_rx_tx_txd),                          //                    .export
		.irq           (irq_mapper_receiver4_irq)                   //                 irq.irq
	);

	Qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c2_clk                                            (altpll_0_c2_clk),                                                    //                                          altpll_0_c2.clk
		.clk_50_clk_clk                                             (clk_clk),                                                            //                                           clk_50_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                 // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                                 //               nios2_gen2_reset_reset_bridge_in_reset.reset
		.TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                     //     TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                             (nios2_gen2_data_master_address),                                     //                               nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                         (nios2_gen2_data_master_waitrequest),                                 //                                                     .waitrequest
		.nios2_gen2_data_master_byteenable                          (nios2_gen2_data_master_byteenable),                                  //                                                     .byteenable
		.nios2_gen2_data_master_read                                (nios2_gen2_data_master_read),                                        //                                                     .read
		.nios2_gen2_data_master_readdata                            (nios2_gen2_data_master_readdata),                                    //                                                     .readdata
		.nios2_gen2_data_master_readdatavalid                       (nios2_gen2_data_master_readdatavalid),                               //                                                     .readdatavalid
		.nios2_gen2_data_master_write                               (nios2_gen2_data_master_write),                                       //                                                     .write
		.nios2_gen2_data_master_writedata                           (nios2_gen2_data_master_writedata),                                   //                                                     .writedata
		.nios2_gen2_data_master_debugaccess                         (nios2_gen2_data_master_debugaccess),                                 //                                                     .debugaccess
		.nios2_gen2_instruction_master_address                      (nios2_gen2_instruction_master_address),                              //                        nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                  (nios2_gen2_instruction_master_waitrequest),                          //                                                     .waitrequest
		.nios2_gen2_instruction_master_read                         (nios2_gen2_instruction_master_read),                                 //                                                     .read
		.nios2_gen2_instruction_master_readdata                     (nios2_gen2_instruction_master_readdata),                             //                                                     .readdata
		.nios2_gen2_instruction_master_readdatavalid                (nios2_gen2_instruction_master_readdatavalid),                        //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                       //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                         //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                          //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                      //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                     //                                                     .writedata
		.EEE_IMGPROC_0_s1_address                                   (mm_interconnect_0_eee_imgproc_0_s1_address),                         //                                     EEE_IMGPROC_0_s1.address
		.EEE_IMGPROC_0_s1_write                                     (mm_interconnect_0_eee_imgproc_0_s1_write),                           //                                                     .write
		.EEE_IMGPROC_0_s1_read                                      (mm_interconnect_0_eee_imgproc_0_s1_read),                            //                                                     .read
		.EEE_IMGPROC_0_s1_readdata                                  (mm_interconnect_0_eee_imgproc_0_s1_readdata),                        //                                                     .readdata
		.EEE_IMGPROC_0_s1_writedata                                 (mm_interconnect_0_eee_imgproc_0_s1_writedata),                       //                                                     .writedata
		.EEE_IMGPROC_0_s1_chipselect                                (mm_interconnect_0_eee_imgproc_0_s1_chipselect),                      //                                                     .chipselect
		.i2c_opencores_camera_avalon_slave_0_address                (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),      //                  i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write                  (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),        //                                                     .write
		.i2c_opencores_camera_avalon_slave_0_readdata               (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),     //                                                     .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata              (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),    //                                                     .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest            (~mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                                                     .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect             (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),   //                                                     .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address                  (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),        //                    i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                    (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),          //                                                     .write
		.i2c_opencores_mipi_avalon_slave_0_readdata                 (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),       //                                                     .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata                (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),      //                                                     .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest              (~mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest),   //                                                     .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect               (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),     //                                                     .chipselect
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                                     .chipselect
		.key_s1_address                                             (mm_interconnect_0_key_s1_address),                                   //                                               key_s1.address
		.key_s1_readdata                                            (mm_interconnect_0_key_s1_readdata),                                  //                                                     .readdata
		.led_s1_address                                             (mm_interconnect_0_led_s1_address),                                   //                                               led_s1.address
		.led_s1_write                                               (mm_interconnect_0_led_s1_write),                                     //                                                     .write
		.led_s1_readdata                                            (mm_interconnect_0_led_s1_readdata),                                  //                                                     .readdata
		.led_s1_writedata                                           (mm_interconnect_0_led_s1_writedata),                                 //                                                     .writedata
		.led_s1_chipselect                                          (mm_interconnect_0_led_s1_chipselect),                                //                                                     .chipselect
		.mipi_pwdn_n_s1_address                                     (mm_interconnect_0_mipi_pwdn_n_s1_address),                           //                                       mipi_pwdn_n_s1.address
		.mipi_pwdn_n_s1_write                                       (mm_interconnect_0_mipi_pwdn_n_s1_write),                             //                                                     .write
		.mipi_pwdn_n_s1_readdata                                    (mm_interconnect_0_mipi_pwdn_n_s1_readdata),                          //                                                     .readdata
		.mipi_pwdn_n_s1_writedata                                   (mm_interconnect_0_mipi_pwdn_n_s1_writedata),                         //                                                     .writedata
		.mipi_pwdn_n_s1_chipselect                                  (mm_interconnect_0_mipi_pwdn_n_s1_chipselect),                        //                                                     .chipselect
		.mipi_reset_n_s1_address                                    (mm_interconnect_0_mipi_reset_n_s1_address),                          //                                      mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                      (mm_interconnect_0_mipi_reset_n_s1_write),                            //                                                     .write
		.mipi_reset_n_s1_readdata                                   (mm_interconnect_0_mipi_reset_n_s1_readdata),                         //                                                     .readdata
		.mipi_reset_n_s1_writedata                                  (mm_interconnect_0_mipi_reset_n_s1_writedata),                        //                                                     .writedata
		.mipi_reset_n_s1_chipselect                                 (mm_interconnect_0_mipi_reset_n_s1_chipselect),                       //                                                     .chipselect
		.nios2_gen2_debug_mem_slave_address                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),               //                           nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                           (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),                 //                                                     .write
		.nios2_gen2_debug_mem_slave_read                            (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),                  //                                                     .read
		.nios2_gen2_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),              //                                                     .readdata
		.nios2_gen2_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),             //                                                     .writedata
		.nios2_gen2_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),            //                                                     .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),           //                                                     .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),           //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                      //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                        //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                     //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                    //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                   //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                   //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                        //                                                     .clken
		.sw_s1_address                                              (mm_interconnect_0_sw_s1_address),                                    //                                                sw_s1.address
		.sw_s1_readdata                                             (mm_interconnect_0_sw_s1_readdata),                                   //                                                     .readdata
		.sysid_qsys_control_slave_address                           (mm_interconnect_0_sysid_qsys_control_slave_address),                 //                             sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_control_slave_readdata),                //                                                     .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_address                       (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),             //                         TERASIC_AUTO_FOCUS_0_mm_ctrl.address
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_write                         (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),               //                                                     .write
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_read                          (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),                //                                                     .read
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata                      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),            //                                                     .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata                     (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),           //                                                     .writedata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect                    (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect),          //                                                     .chipselect
		.timer_s1_address                                           (mm_interconnect_0_timer_s1_address),                                 //                                             timer_s1.address
		.timer_s1_write                                             (mm_interconnect_0_timer_s1_write),                                   //                                                     .write
		.timer_s1_readdata                                          (mm_interconnect_0_timer_s1_readdata),                                //                                                     .readdata
		.timer_s1_writedata                                         (mm_interconnect_0_timer_s1_writedata),                               //                                                     .writedata
		.timer_s1_chipselect                                        (mm_interconnect_0_timer_s1_chipselect),                              //                                                     .chipselect
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                                //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                                  //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                                   //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                               //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                              //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                          //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                              //                                                     .chipselect
	);

	Qsys_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c2_clk                                 (altpll_0_c2_clk),                          //                               altpll_0_c2.clk
		.alt_vip_vfb_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // alt_vip_vfb_0_reset_reset_bridge_in_reset.reset
		.alt_vip_vfb_0_read_master_address               (alt_vip_vfb_0_read_master_address),        //                 alt_vip_vfb_0_read_master.address
		.alt_vip_vfb_0_read_master_waitrequest           (alt_vip_vfb_0_read_master_waitrequest),    //                                          .waitrequest
		.alt_vip_vfb_0_read_master_burstcount            (alt_vip_vfb_0_read_master_burstcount),     //                                          .burstcount
		.alt_vip_vfb_0_read_master_read                  (alt_vip_vfb_0_read_master_read),           //                                          .read
		.alt_vip_vfb_0_read_master_readdata              (alt_vip_vfb_0_read_master_readdata),       //                                          .readdata
		.alt_vip_vfb_0_read_master_readdatavalid         (alt_vip_vfb_0_read_master_readdatavalid),  //                                          .readdatavalid
		.alt_vip_vfb_0_write_master_address              (alt_vip_vfb_0_write_master_address),       //                alt_vip_vfb_0_write_master.address
		.alt_vip_vfb_0_write_master_waitrequest          (alt_vip_vfb_0_write_master_waitrequest),   //                                          .waitrequest
		.alt_vip_vfb_0_write_master_burstcount           (alt_vip_vfb_0_write_master_burstcount),    //                                          .burstcount
		.alt_vip_vfb_0_write_master_write                (alt_vip_vfb_0_write_master_write),         //                                          .write
		.alt_vip_vfb_0_write_master_writedata            (alt_vip_vfb_0_write_master_writedata),     //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_1_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_1_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_1_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_1_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_1_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_1_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_1_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_1_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_1_sdram_s1_chipselect)     //                                          .chipselect
	);

	Qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c2_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
